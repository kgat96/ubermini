* F:\appotech\opcode\ubertoothp\hardware\t1.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/11/2016 13:13:09

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  Net-_C1-Pad1_ Net-_C1-Pad2_ R		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ CP		

.end
